x1 x2 x3 x4 x5 
0.7951248 1.4659937 0.8494663 -0.495743 1.1296365 
0.6492540 0.4383383 -0.082964 -0.159053 0.3414969 
0.3293332 -0.195318 0.0923112 -0.398622 -0.029444 
-0.288707 0.9564703 1.3740610 -1.338867 1.0681129 
-0.274006 -0.660734 -0.649236 0.4974154 -0.382859 
0.8689484 1.6575051 1.5991888 -1.159828 1.6806745 
-0.162992 -0.995362 -1.209802 0.8596714 -0.924777 
-0.587805 -0.537352 0.1345542 0.8285142 -0.387999 
-0.657559 -0.587003 -0.221320 -0.906280 -0.484596 
-0.601995 0.1742395 0.8128345 -0.250058 0.1806672 
-0.405701 0.7508328 1.6372188 -0.406460 0.8170545 
0.8720166 1.2059380 0.4706571 0.6126053 1.1016069 
0.7753430 1.6083786 1.3338184 -0.344012 1.0746955 
-0.788343 -1.759760 -1.216673 1.8386653 -1.659841 
-0.593654 -0.041819 0.2437219 0.5314528 -0.168301 
0.3001320 -0.067325 -0.065440 0.6050985 -0.320503 
-0.065989 -0.517402 -1.073068 0.2219711 -0.681583 
-0.319732 -0.648886 -0.146921 0.4182412 -0.600338 
-0.300885 -0.954441 -1.780613 0.7245473 -0.987820 
0.9765962 1.5668784 0.4230049 -0.823279 1.4826839 
0.4307993 0.6454005 0.8938824 -1.390935 0.7291835 
-0.966377 -2.317104 -1.429936 0.8993891 -1.748596 
-0.085559 -0.613411 -0.253470 0.2577651 -0.585119 
-0.117789 0.8263267 1.1811796 -0.957771 0.6881731 
0.0344681 -0.636843 -0.855790 0.8868225 -0.606171 
-0.090756 -0.087809 0.2127512 -0.923705 -0.067943 
-0.401492 -0.641932 -0.907291 0.9523962 -0.788080 
0.1194116 0.1167911 -0.841477 0.6790472 0.0192483 
-0.062365 0.1333660 -0.064575 0.0470881 0.2125302 
0.3867436 0.8669972 0.5507640 -1.193653 0.8720201 
0.8026807 0.8528774 0.3209627 -0.802955 0.9530817 
-0.179739 -0.117645 -0.053033 -0.470771 -0.089321 
0.5324187 1.6661851 1.8500792 -1.511553 1.6616919 
-0.703566 0.1383046 0.7942693 -0.783776 0.4346688 
-0.286153 -0.938862 -1.646141 0.3122314 -0.709328 
0.1131143 0.7729262 0.4243400 -0.591867 0.6212415 
-0.783578 -0.366132 0.2969030 -0.716619 -0.519068 
0.5692348 -0.046606 -0.462934 0.4809312 0.0058366 
0.0644239 0.0292505 0.1107860 -0.229817 -0.070709 
-0.385989 -0.259179 -0.435270 -0.208291 -0.198529 
0.4640754 0.1685348 -0.178911 -0.084619 0.3700194 
0.4459827 1.9335389 2.4455264 -1.475687 2.0414369 
0.6162926 0.2465663 -0.368012 -0.095003 0.0418567 
-0.156246 -0.099045 0.4662705 0.7290251 -0.182159 
0.8091675 0.4165856 -0.774343 0.5823631 0.4286500 
-0.760782 -0.841854 0.7824814 1.1208487 -0.917386 
0.0098548 -0.251564 -0.392787 -0.664964 -0.227211 
-0.828865 -1.048615 -0.532274 0.3896414 -1.138607 
0.1541587 -0.709360 -2.388692 0.7633626 -1.040224 
0.2061637 -0.059131 -1.378504 0.1628405 -0.013058 
0.2863743 0.3104169 0.6985656 -1.400817 0.3513958 
0.6292003 0.4616197 0.2776306 -0.175387 0.2528633 
0.6746381 -0.569481 -1.548959 0.3730588 -0.533666 
-0.750104 -1.893544 -1.930970 1.0350515 -1.625937 
0.6427851 1.1493254 0.9881173 -1.206013 1.4705501 
0.8533874 1.1251147 1.4291152 -1.121772 1.3759816 
-0.643284 -0.801159 -0.963902 -0.351585 -0.854083 
0.4712938 0.1966518 0.0983572 0.4922122 0.4015961 
-0.467282 0.0936705 1.1333452 0.5846135 0.0767836 
0.0041952 -0.440372 -0.815910 0.4366609 -0.297846 
0.9406344 1.7505747 0.3554521 -2.556127 1.9048797 
-0.217721 0.6154592 0.9060832 -1.009213 0.8392086 
-0.256243 -1.466090 -2.127546 1.0557487 -1.184909 
-0.340582 -0.356630 0.1227193 0.6423055 -0.246373 
-0.026168 -0.320818 -0.509866 0.3917304 -0.116677 
-0.615064 -0.209531 -0.520082 -0.951801 -0.217512 
-0.819663 -0.983347 0.0735845 1.5540028 -0.824734 
0.8288736 0.8039635 -0.373348 -0.444381 0.8669299 
-0.747015 -0.665767 0.4149621 1.3871703 -0.517551 
0.9667007 2.4353076 1.5362534 -2.052017 2.1172288 
-0.845485 -1.256079 -0.556444 0.2315288 -1.439777 
-0.374029 -1.125133 -1.317344 2.2365211 -0.979354 
-0.898795 -0.687607 0.6009825 0.7682289 -0.377159 
0.8944059 1.5772605 0.8852084 -1.076970 1.5929353 
0.6479262 0.6607607 0.5361878 0.3522877 0.8848895 
-0.611293 -1.210511 -0.859292 1.2482944 -1.162151 
0.3352886 -0.581449 -0.945076 0.6830510 -0.454137 
0.4609838 0.5409692 -0.309208 -0.204082 0.4600558 
-0.651810 -0.884146 -0.537106 0.1188759 -0.818837 
0.6251817 0.2499355 -0.079492 0.0107955 0.2361106 
-0.938598 -0.863434 -0.155008 0.6282431 -1.063052 
-0.606190 -0.322794 -0.527588 0.0575769 -0.637832 
-0.696893 -1.742968 -2.212388 1.7213980 -2.138510 
0.9707394 2.9338285 2.2716376 -1.991643 2.7324361 
-0.362486 -1.433526 -1.863661 1.6354141 -1.189069 
0.3421594 -0.158149 -0.396428 0.0211211 -0.401455 
-0.308264 -0.875173 -1.677259 0.8759929 -0.889976 
0.5887926 1.3614914 1.3065834 -1.272100 1.2413254 
-0.890234 -0.924308 -0.468239 1.2736622 -1.294625 
-0.202667 -0.286784 0.3981495 0.4245548 -0.009541 
-0.409286 -0.063299 0.3260226 0.0726959 -0.127146 
0.0891216 -0.429723 -1.002515 0.5297188 -0.432764 
0.4974958 0.7377782 -0.292009 -0.194963 0.4535805 
0.9845518 2.6705953 2.7554433 -2.142764 2.5642140 
-0.472496 0.2559677 0.9359239 -0.721113 0.2873916 
0.2520343 -0.722629 -0.947907 1.2661002 -0.656331 
-0.476973 0.9294276 1.9026163 -1.954383 1.1187862 
-0.320654 -1.271623 -1.567543 0.6498468 -1.116025 
-0.633306 -0.512073 -0.091336 0.4624494 -0.370662 
-0.848356 -1.319060 -0.339990 0.6918319 -0.896382 
-0.181378 -0.404727 0.1071440 1.0646224 -0.268156 
0.5077253 0.7279662 0.0537159 -1.263132 0.5359427 
0.1637997 -0.007619 -0.410745 -0.746450 -0.058405 
0.4879797 0.8903853 0.8273497 -0.295608 0.4920035 
-0.908983 -1.675592 -0.553373 0.9668363 -1.758852 
-0.103566 -0.398673 0.1978061 0.3812289 -0.180530 
0.3808031 -0.109223 -0.723062 0.3582780 0.0623570 
-0.729576 -0.294755 -0.877098 -0.608904 -0.395139 
0.6969510 0.7202851 0.3863920 0.0017413 0.6675553 
-0.437015 -1.024901 -1.409996 0.1841990 -1.095813 
-0.616184 -0.280946 0.2284848 0.2467084 -0.150116 
-0.733658 -1.081059 -0.495434 0.2970100 -1.117277 
0.7705527 0.6756519 -0.130704 0.5023930 0.7662096 
-0.995054 -2.121065 -0.893041 0.7883965 -1.519340 
-0.912628 -1.147811 -1.028005 0.7403726 -1.380872 
0.3460033 -0.052989 -0.321623 -0.065574 0.1612174 
-0.709059 -0.714296 -0.008790 0.6955404 -0.743896 
-0.128492 0.5574071 1.1376622 -0.629407 0.7616965 
-0.798517 -1.664436 -0.868440 1.1134115 -1.925653 
0.6092068 -0.622198 -1.258502 0.8513871 -0.327293 
0.6606706 0.9900374 0.3381230 -0.683266 0.9554618 
-0.277440 -0.136806 0.7372290 0.9085125 -0.231344 
0.2907204 0.3691711 0.1583181 -0.086507 0.5036044 
0.5617941 0.3486212 0.0488140 -0.117754 0.3322341 
-0.313722 -0.189013 -0.024487 -0.322503 -0.352531 
-0.860993 -0.015281 0.3314121 -0.362565 -0.270424 
-0.589587 -0.407711 0.1411205 0.7147475 -0.132899 
-0.547547 -0.744390 -0.404346 0.2909553 -0.647048 
0.2405824 1.9046074 3.8120837 -1.744249 1.7703864 
0.4202369 0.5076182 0.4399383 -0.649645 0.4870985 
0.5640835 0.4014689 -0.769117 -1.364028 0.3892776 
0.7847565 1.4556455 0.5627938 -0.974648 1.2852250 
0.6891642 0.4241370 -0.847041 0.2865062 0.3652687 
-0.359458 -0.849471 -0.935474 1.3099703 -1.082647 
-0.498425 0.5469988 1.1076139 -0.988642 0.6687146 
-0.944079 -0.992920 -0.114031 0.8377348 -1.013309 
-0.940151 -1.822900 -1.014141 0.8692064 -1.410962 
-0.707131 -2.062312 -1.026705 1.7799789 -2.032058 
-0.961545 -2.447186 -1.728186 0.3465052 -2.283678 
-0.264836 -0.533567 -0.033540 -0.263758 -0.342911 
0.8622754 1.9996237 2.1406665 -1.605749 2.1995827 
-0.055747 -1.168291 -2.037211 0.7806095 -1.131721 
0.2814351 -0.127743 -0.568576 1.2972471 -0.293990 
-0.413613 0.1423629 0.2941597 -0.235570 0.1229056 
0.8907116 0.9971883 -0.542431 -0.200727 0.6501760 
-0.051131 0.1973085 0.7682554 -0.281564 0.0682150 
0.8188878 1.1917751 1.0601473 -1.086228 1.0837724 
-0.164528 0.3766261 1.5682804 -0.984926 0.6084364 
0.6074776 1.2590114 1.3848319 -1.901943 1.2502649 
-0.254204 0.4545548 0.8911672 -0.329669 0.1579526 
-0.957638 -1.830779 -0.173446 1.4371561 -1.553117 
-0.557921 -0.071999 0.3693986 -0.103176 -0.216655 
-0.480003 -0.706073 -0.244528 0.1577212 -0.511190 
0.3707818 1.2260185 1.5134422 0.0388854 1.1889469 
-0.205712 0.6240025 0.1510036 -0.177369 0.1184109 
0.3379701 0.3386953 -0.124865 -0.074330 0.4738808 
-0.337110 0.2743549 0.3949042 -1.048195 0.2457547 
0.8333700 1.8723020 1.7662108 -1.582851 1.8171326 
-0.779304 -1.111330 -0.786981 1.6978544 -1.316691 
-0.872103 -1.577743 -1.328775 1.3325137 -1.475024 
-0.793598 -1.397824 -1.277083 1.7706498 -1.287261 
-0.512527 -1.099316 -1.188200 0.7333407 -1.526522 
0.8993936 1.6009769 1.1213339 -0.423348 1.7452875 
0.7228831 0.8188044 0.3673160 0.4028884 1.0049467 
0.9197444 1.7033989 0.6851569 -0.918919 1.7016325 
0.1796201 -0.763431 -1.723474 1.3197080 -0.675046 
0.4769924 0.4056957 -0.441877 0.1755571 0.3249506 
-0.539636 0.5480275 1.0923351 -0.837386 0.7892780 
0.0129175 -0.437565 -0.431557 -0.382268 -0.434563 
0.3115237 0.7126962 1.2249449 -0.962805 0.7545177 
0.3960875 0.0672630 0.8486665 -0.731294 0.4325944 
0.1473792 -0.421800 0.2546549 1.5684284 -0.472511 
-0.758090 -1.642334 -1.316013 0.3224856 -1.477563 
-0.622916 -1.136036 -0.705720 1.0268277 -1.074525 
-0.268431 -0.083632 0.3074316 0.5727216 -0.407180 
-0.719888 -1.010353 -1.233676 0.4102866 -1.256121 
0.9468853 1.2941902 0.4557417 -1.447969 1.3869945 
0.5433529 1.0237692 0.9470995 -1.027045 1.1703737 
-0.071841 0.5157852 0.7277789 0.0408175 0.5674031 
0.2717747 0.0342518 0.4387345 -0.051832 0.0842485 
-0.916801 -1.873547 -0.515568 1.9448677 -1.889474 
0.4188064 0.8569235 1.0717841 -0.637271 0.3134675 
-0.208381 -0.669963 -0.574304 0.7068947 -0.590488 
-0.378870 -1.389977 -1.383351 1.0522604 -1.101952 
-0.838937 -0.861449 -0.106238 -0.014886 -0.935757 
0.3150792 -0.680414 -0.961002 1.1383428 -0.731317 
-0.902786 -1.330934 -0.929778 1.3554989 -1.457280 
0.4759289 0.4972126 0.4970745 -0.466469 0.5879626 
-0.299477 0.5039738 1.2974600 -1.678713 0.5610453 
-0.448530 -2.050997 -2.071915 2.3325184 -1.828659 
0.9117133 1.7171028 1.3918468 -1.036501 1.9258757 
-0.880494 -2.648205 -2.293240 2.0944258 -2.735627 
-0.754338 -1.690675 -1.575753 1.4804020 -1.577183 
0.7523936 0.3901343 0.1035568 1.2155767 0.6304247 
-0.738024 -0.603746 -0.141822 0.5506758 -0.614872 
-0.038442 -0.425802 0.3132979 0.5977404 -0.278165 
0.1489239 -0.911429 -1.642520 0.5188925 -0.865078 
-0.996101 -2.175634 -0.563014 2.2829132 -2.206809 
-0.155241 -0.557258 -0.315784 0.2049723 -0.529314 
-0.139696 0.3567063 1.2466315 0.4757922 0.5126378 
0.5002685 -0.035274 -1.291757 0.0985165 -0.304267 
-0.787908 -1.481539 -1.042425 1.3675652 -1.820967 
0.6793598 0.4955353 0.4583944 0.0778570 0.6761310 
0.2944486 0.4672015 -0.018304 -1.560487 0.5176180 
0.1250385 0.2146189 0.2525907 -0.292297 -0.152957 
-0.429911 0.9318860 1.7802884 -1.195618 0.7182710 
0.7172907 1.2397591 0.9122603 -0.244591 1.0496295 
-0.188193 -0.748281 -0.300827 1.0734840 -0.748703 
-0.230042 -0.387344 -0.271749 0.3161172 -0.543824 
0.2360750 -0.494915 -1.433972 -0.078507 -0.578011 
0.5743075 0.5769022 0.2719260 0.1933730 0.6407329 
0.2510495 0.0538576 0.0129357 0.1282797 0.3953071 
0.9743992 2.0193709 1.9870513 -0.688308 1.9797549 
0.4266830 0.9506305 1.6107041 -1.414112 1.3448499 
-0.185593 -1.551133 -1.906497 2.4471486 -1.975031 
-0.510131 -1.409885 -1.402729 0.5164282 -1.604471 
0.0184213 1.4854883 2.1444638 -2.908319 1.4531811 
-0.226279 0.2309864 0.3347362 0.3594566 -0.260622 
0.4087878 -0.766586 -1.488972 0.8817696 -0.697276 
-0.468018 -0.686676 -0.596158 0.7517812 -0.537722 
-0.369964 -0.224398 0.5977939 0.8437741 -0.207746 
0.5175655 1.1758609 1.6600837 -0.842866 1.1096460 
-0.768170 -2.818203 -2.559008 1.6663901 -2.633709 
0.2009710 0.2668262 0.0613525 -0.479911 0.6035055 
-0.033655 -0.337766 -0.605390 -0.185898 -0.017856 
-0.240210 -0.011341 0.9843497 -0.394991 0.1448789 
0.6956779 1.7913906 1.8701811 -1.252052 1.8376761 
-0.282702 0.0765031 1.2072621 1.0981696 -0.171591 
0.2757441 -0.783673 -1.970982 0.9954999 -0.836243 
-0.017310 -0.599000 -0.653011 0.4145143 -0.549470 
-0.244014 -0.496485 -0.193985 0.5100745 -0.621281 
0.3903312 1.6299365 2.2412625 -1.929283 1.3386098 
0.0943508 0.6630182 0.4833398 -1.504326 0.6355177 
-0.671992 -1.014502 -1.062826 0.6146287 -1.242405 
-0.047274 0.5706305 0.6201884 -0.147070 0.5802384 
-0.626516 -0.815802 -0.449909 1.8896667 -0.803906 
0.9974337 2.1762300 0.5780095 -1.130419 1.9465076 
-0.149042 0.0086390 0.1393206 0.2509225 -0.160116 
0.0806680 -0.219573 -0.891628 -0.538828 0.1885994 
-0.001712 0.8969091 0.7907430 -0.554005 0.9225565 
-0.721791 -0.888786 -1.008516 0.0182684 -0.796680 
0.9572578 0.8717234 -0.012631 -0.708030 1.1648178 
-0.532994 0.1302695 0.2871983 -0.254874 -0.444231 
0.4159178 -0.175662 -0.489906 0.1554081 -0.341654 
-0.922250 -2.403060 -2.776067 1.1347818 -2.368113 
-0.030797 0.0608981 0.1635075 0.9909198 -0.139894 
0.1118505 0.3846037 0.7006467 -0.437729 0.2183842 
0.3220207 1.1659782 1.4500187 -1.690305 1.1363015 
-0.815348 -1.605760 -0.757901 2.1811120 -1.221646 
0.1227273 -0.344038 -0.164006 0.1484418 -0.358284 
0.9508609 1.9564282 1.1106746 -1.843687 2.1915807 
-0.367915 -0.466370 0.0321735 -0.038594 -0.321447 
0.3604824 0.3346543 0.6593682 -0.218769 0.7240746 
0.3578073 1.0696099 1.5409477 -0.528787 1.4465131 
-0.855303 -1.930604 -1.515041 2.7413325 -2.417656 
-0.235278 -0.101740 -0.199708 -0.452191 0.0528633 
-0.304749 0.1567538 1.7457775 -0.059661 0.4145030 
0.2251026 0.0445069 -0.264884 0.7029901 -0.109294 
0.7994640 1.7579965 1.1533690 -1.227980 1.5392502 
-0.953438 -1.181908 -0.240353 0.6666060 -1.352739 
0.0462404 0.6836122 1.4091859 -0.678817 0.3629437 
0.3165954 0.7522574 0.5173745 -1.352236 0.4478258 
-0.487537 -0.840202 -0.613063 0.4714603 -0.881470 
-0.121078 0.1064109 0.0093285 -0.006858 0.0483033 
0.4027071 1.0459404 1.5051024 -0.417245 1.0330877 
-0.821147 0.0370016 1.1711563 -0.936645 0.1288716 
0.8071501 1.3811369 0.6331886 -1.813774 1.4239022 
-0.766928 -0.787325 0.2120515 1.4049884 -0.776494 
0.9077734 0.3943878 -0.686108 0.1431584 0.2602402 
-0.834270 -0.733019 -0.261431 0.8143907 -0.811819 
0.3759794 1.2694710 1.2879803 -1.136201 1.0397709 
0.1747322 0.5999288 0.1888732 -0.308972 0.5988400 
0.2584634 0.4094523 -0.185286 0.2101630 0.2693813 
0.7422560 1.0161588 0.7438244 -1.033940 1.0893789 
-0.561336 -0.149439 0.9956963 -0.141179 0.1695144 
0.5381312 -0.205523 -0.480723 0.6331393 -0.250885 
-0.712949 -0.078033 0.0225373 0.0268391 -0.188517 
0.4489263 0.7634920 1.2488553 0.1351947 0.7334327 
0.7507519 1.0910281 0.9218679 -1.168875 0.9957364 
-0.394616 -0.483857 -0.811911 0.5443870 -0.908450 
0.1336779 -0.384287 0.0698417 0.1988312 -0.121024 
0.2978572 0.8806458 0.8139681 -0.795772 0.8094807 
0.0264832 0.8306883 0.6109642 -0.771746 0.7051804 
-0.680505 -1.372522 -1.265228 -0.369685 -1.202971 
0.9249691 1.5272208 0.1936551 -0.871588 1.2070636 
0.8277898 1.0094248 0.6733235 -0.270205 1.2192130 
0.5941359 -0.179024 -0.344039 0.5705211 -0.052414 
0.7116145 1.2316063 1.4660094 -1.055056 1.5702775 
-0.527762 0.0172631 0.5228033 -0.489982 0.1046983 
-0.576329 0.2245320 0.5274747 -0.861787 0.1136093 
-0.133923 -0.655491 0.0173395 0.4462451 -0.474893 
0.4067701 -0.348659 -0.379960 0.9012549 -0.284870 
-0.581729 0.3044766 -0.104314 -1.751786 0.4192745 
-0.011963 0.5196487 0.3611175 -0.375404 0.6144511 
-0.391257 0.9435577 1.6994688 -0.887646 1.2284275 
0.5096140 -0.362335 -0.918323 0.1235897 -0.196061 
0.3275741 0.2800474 -0.830384 -0.734343 0.4962283 
0.1673214 0.3218409 0.5727461 -1.428530 0.5471320 
0.5140757 0.9077635 1.1636850 -0.942517 0.9104196 
0.8152549 0.3453964 -0.804699 -0.063994 0.5584955 
-0.462278 -0.547686 -0.675922 0.9605708 -0.416186 
0.8363724 1.8098453 1.8053515 -2.824486 1.7080686 
-0.858768 -1.531760 -1.838938 1.1465606 -1.852954 
0.9606723 2.1024375 1.7166014 -1.437335 2.3194622 
-0.348913 -0.165174 -0.166535 -1.092846 -0.080804 
-0.333722 -0.461417 -0.477010 -0.700640 -0.610726 
0.8491436 0.5595540 -1.126161 0.3414332 0.1516593 
0.9543080 1.3513917 0.9780966 -0.696249 1.4931587 
-0.678658 -0.970507 0.1200952 0.5578364 -0.734083 
0.6674682 0.0995424 -0.378652 -0.313765 0.2534373 
-0.725928 -2.246431 -2.487727 2.1075137 -2.158883 
0.9224380 2.3195851 2.3812885 -2.286092 2.3424523 
-0.456990 -0.503639 -0.673099 0.3351284 -0.571472 
0.0316823 0.2952087 0.5911926 0.4292895 0.3209545 
0.0745893 -0.468308 -0.608365 0.9811801 -0.654469 
0.6207564 0.1866514 -0.460277 0.0651278 0.4424648 
0.9032662 2.5993027 2.5871150 -2.377643 2.8968862 
0.7020434 1.4225303 1.1908073 -1.247737 1.2027396 
-0.221841 -1.067508 -0.877949 1.4297824 -0.952796 
0.7132210 0.1229917 -0.692748 0.3280118 0.0223367 
0.4913584 -0.244627 -0.578585 0.2770081 -0.102704 
0.6586732 0.3285609 -0.287954 0.1139228 0.2410986 
-0.195904 0.0872228 -0.350753 -0.619456 -0.306481 
-0.549255 -0.901504 -1.200362 1.0149279 -1.336807 
-0.174274 -0.302153 0.8009630 -1.002397 -0.035377 
0.0791080 -0.032262 0.1271493 0.1053676 -0.164737 
-0.692531 -0.778546 0.0801579 0.3642345 -0.831587 
0.1903928 -0.562176 -1.058801 0.9769749 -0.467056 
-0.012332 -0.029044 0.4316074 1.4672090 -0.280273 
-0.978359 -1.563819 -0.025555 1.5809582 -2.003516 
0.9950465 1.2871509 0.2026086 -0.288389 1.4024792 
-0.555199 -1.351036 -0.747626 1.1849433 -0.871565 
-0.124795 -0.115304 -0.043671 -0.512371 0.0370798 
0.1960787 -0.182511 -0.825474 0.2383770 0.0294265 
-0.023074 0.4179295 0.6147301 -0.340307 0.4718328 
0.0221349 0.5337485 0.1702386 -0.603233 0.4113746 
-0.445315 -0.699562 -0.189941 1.5235308 -0.857578 
-0.647983 -0.833561 -1.084485 -0.121308 -0.760937 
-0.691752 -1.284963 -0.663606 1.8184662 -1.700778 
0.0602407 -0.729350 -1.505545 1.2378954 -0.479873 
-0.099706 -0.946985 -1.815701 1.5903575 -0.771955 
-0.500160 0.1824872 0.0555999 -0.426032 0.0588004 
-0.327545 -0.484687 -0.425825 0.8007867 -0.425146 
0.5564478 1.3272933 1.9389170 -1.478265 1.6085620 
0.0545391 0.2338000 -0.087477 -1.100002 0.3036718 
-0.424200 -0.152776 0.9277851 -0.335633 -0.143295 
0.0414940 0.1658038 0.7770295 -0.132661 0.3799175 
-0.095057 -0.796996 -1.181713 1.2263540 -0.692043 
-0.879047 -0.314782 0.4891854 -0.647685 -0.046290 
-0.986002 -1.609221 -0.156155 1.7411281 -1.394646 
-0.904482 -3.033997 -3.131589 3.1880503 -3.088466 
0.1842666 0.2024597 0.4123610 -0.671014 0.2089399 
0.7596959 0.9814348 0.0891330 -1.715528 0.8534860 
0.9380058 0.9771879 0.6511407 -0.568554 1.0564828 
0.6124119 1.1097273 0.7235095 -1.301101 0.7722006 
0.2666370 -0.414374 -0.783218 0.0060843 -0.114241 
0.9349986 1.3746248 0.8684541 -0.222870 1.4117113 
-0.432377 -0.379274 0.5423324 0.3084556 -0.631048 
0.9901400 2.3575888 1.3279883 -1.652418 2.4670624 
0.0980834 1.0295653 0.8575410 -0.833728 1.1824268 
-0.800689 -1.710483 -1.698032 1.6212333 -1.504431 
-0.572592 0.1111910 1.0698023 -0.025545 0.1056177 
0.5258095 1.1432269 1.195373 -0.586478 0.9231320 
0.7804052 1.3326398 0.7141924 -0.450623 1.3095146 
0.8811221 1.0989298 -0.728811 -0.896899 1.1485841 
0.4361229 -0.369922 -1.157743 0.5893927 -0.359818 
0.0507959 -0.454438 -0.585708 0.2616278 -0.045017 
0.0861597 0.0149408 -0.298150 0.6467931 -0.002215 
0.0031157 0.9656732 0.6253770 -1.066788 0.9353577 
-0.168439 0.4696610 0.0813883 -0.127370 0.1471291 
0.9318597 0.1009498 -0.333934 1.4149072 0.0332738 
-0.639774 -1.515249 -1.353568 1.1728308 -1.229740 
0.1419538 0.6940108 0.1727312 -1.374985 0.5715168 
0.4577745 1.5122711 1.0846819 -2.222079 1.5093449 
0.7379023 0.9222034 0.5844278 0.1706369 0.8276281 
-0.674738 0.1468339 0.9458019 0.2727073 0.2934448 
-0.741113 -1.306410 -1.604720 0.9319159 -1.608001 
-0.196362 -0.257256 -0.657932 -0.108287 -0.554005 
0.8579695 1.8309779 2.0639212 -1.317141 1.8775075 
0.0565639 0.4777311 0.5654774 -0.636760 0.2793166 
-0.249123 0.2740095 1.0057102 -0.523045 0.3104503 
-0.260194 -0.296627 -0.205325 -0.532399 -0.336807 
-0.529989 -0.573362 0.5357787 0.3972114 -0.559660 
-0.115036 0.6506206 0.5584011 -1.307590 0.6604650 
0.9833102 2.2391879 0.4922795 -1.634112 1.7979963 
0.7623733 0.6092540 -0.360250 1.1008076 0.3457494 
-0.654167 -1.236816 -1.170794 0.8089882 -1.422768 
-0.772334 -0.331132 0.2204853 0.2268119 -0.634453 
-0.144376 -0.230180 -0.236701 -0.597212 -0.369111 
-0.970446 -1.991968 -1.151024 1.1885538 -1.556582 
-0.930570 -1.220047 -0.251982 1.1558019 -1.150913 
0.6550090 0.5868974 -0.716950 0.0685881 0.1311248 
0.2165496 0.4834243 0.2844063 -1.220202 0.5347567 
0.5786582 0.5299625 0.2232585 -0.238167 0.9064594 
-0.516906 0.4467629 1.2608437 -0.153043 0.3980999 
0.6393757 1.2052306 1.5805743 -0.758657 1.0117528 
0.5977398 0.3130729 -0.451548 0.1058377 0.3570603 
0.7316541 0.7431713 0.6891327 -0.023067 0.2681420 
0.4411741 0.5913934 0.6675324 0.3749913 0.8884900 
0.8641401 1.5517867 0.7467211 -1.787707 1.5300956 
0.7269876 0.7703907 -0.276727 0.1867246 0.6478209 
-0.599490 -0.235480 0.7551978 0.0828448 -0.492779 
0.8845085 0.9115765 0.2636508 -0.618716 0.9940823 
0.5288500 0.0582256 -1.093124 1.3412333 0.0126578 
0.1825045 0.6382539 0.6473407 -0.317021 0.7432050 
-0.419203 -1.295561 -1.529494 1.9172879 -1.270066 
0.1568188 -0.395417 -0.035844 2.0074473 -0.310794 
0.1307790 0.7971669 1.3604316 -0.190943 0.7115253 
0.2224749 -0.022690 0.0298193 -0.461297 0.1822138 
0.6353148 0.8115493 -0.133799 -0.775469 0.8032108 
-0.005668 -0.269943 -0.222533 -0.475007 -0.064668 
0.9151439 2.077667 1.2802071 -2.168255 2.0738022 
-0.453110 -0.332426 -0.628400 -0.433290 -0.457587 
0.2622556 0.1512198 0.2426988 -0.000978 0.5917149 
-0.924134 -1.785563 -1.607339 0.9200628 -1.709897 
0.3948472 1.4378863 1.6680693 -2.488477 1.5845599 
-0.396209 -1.040725 -1.295216 1.4534453 -0.999411 
0.8477927 0.3708589 -0.117522 0.3054047 0.4634967 
0.1923765 0.0727153 -0.059541 -0.810896 0.1972082 
-0.982866 -1.505245 -0.759436 1.0872837 -2.057534 
0.2289049 1.0613702 1.0152487 -0.367112 0.8945081 
0.2781375 -0.919045 -0.707345 0.7970437 -0.907606 
-0.077740 -0.197604 -1.135153 0.2336391 0.0010038 
-0.842552 -0.824185 -0.624472 -0.099726 -0.971552 
0.3537500 0.1796575 0.0443823 -0.031538 0.5512275 
-0.932938 -1.424442 -0.329234 1.1983102 -1.356470 
-0.382529 0.6722160 0.3032524 -0.741865 0.5217743 
0.7777649 1.2714976 0.8377667 -0.883412 1.6313070 
-0.989306 -1.132277 -0.387563 -0.259930 -1.165284 
0.6682720 1.3158620 1.0355633 -1.870774 1.2796554 
0.3665159 -0.478411 -0.913643 0.0938380 -0.448463 
-0.504422 -0.306081 0.2673303 0.5628887 -0.238851 
-0.867809 -0.609098 0.0351099 -0.549999 -0.722055 
0.7068150 1.0731628 0.3429607 -0.789869 1.2939515 
0.5460594 1.0398317 0.9544200 0.0861650 0.6848930 
-0.330610 0.7848364 0.6785461 -0.278709 0.2029613 
0.6815516 0.8448846 0.1856585 -0.762904 0.7474032 
0.7674507 0.4330294 -0.422891 0.4881340 0.1756758 
0.5555414 0.0492190 0.5091399 -0.165162 0.0942214 
0.4837652 0.4861773 0.7606081 -0.660618 0.8615776 
-0.237994 0.2417464 1.4889413 -0.137333 0.2840175 
-0.040628 0.0803126 -0.099960 -0.572957 0.1926457 
0.5210098 0.6298677 1.0452170 0.6577414 0.2252121 
-0.804196 -1.078280 -0.354132 0.9233314 -1.035957 
0.0395674 -0.931910 -1.244024 1.2325293 -0.504793 
0.2320163 0.3631117 0.1490197 -0.356226 0.9400913 
0.4343509 -0.001294 -0.048281 0.4612479 -0.094548 
0.5802748 0.7133363 1.3491055 -0.168286 0.9858594 
-0.109400 -0.094488 0.3819954 -0.855837 0.0964325 
-0.294230 -0.968310 -0.694449 0.2154211 -0.663373 
-0.352207 0.6009587 1.0258552 -0.513165 0.4821808 
-0.495679 -0.807975 -1.449765 0.4527023 -1.019946 
-0.522169 -0.120840 0.4504053 0.0544573 -0.256423 
-0.540945 -0.266602 0.3784200 -1.523420 -0.035075 
-0.423024 -1.062212 -0.503146 1.8803858 -1.208387 
-0.567835 -0.142147 -0.213644 -0.818099 -0.419167 
-0.080127 -0.168254 -1.143449 -0.504187 -0.097426 
0.2101664 1.4054488 1.9604085 -1.544807 1.2658606 
-0.072418 -0.130834 -0.736352 -0.300243 -0.206771 
0.8213769 1.3963007 2.0204064 -0.581888 1.3198758 
-0.628273 -1.093431 -1.048801 0.4440726 -1.367079 
-0.056043 -1.244335 -0.497297 1.5019349 -0.968651 
-0.663778 -0.589417 -0.317860 -0.216093 -0.670211 
0.1367928 -0.213665 -1.098525 -0.050117 -0.233663 
0.5484410 -0.523702 -1.341186 0.7558112 -0.568454 
0.7471076 0.6364994 -0.001549 -0.909970 0.7855112 
-0.811915 -0.752878 -0.592382 0.7754375 -0.843338 
0.3764265 0.2936814 0.4017411 -0.543694 0.2973623 
0.4927599 0.7900383 0.9676406 -0.867565 0.8238275 
-0.687646 -1.959299 -2.175755 2.5627571 -1.776750 
0.6035813 0.8390644 0.2339692 -0.498716 0.9772092 
-0.215231 1.0818684 1.4379305 -2.071580 0.8425354 
-0.666337 -1.204104 -0.413295 0.9448076 -0.942210 
0.0683466 0.2112378 0.8740230 0.8255017 0.2324464 
0.2141114 0.4417738 0.3478639 -0.113283 0.3802713 
-0.892820 -1.450890 -1.111701 1.2869192 -1.677597 
-0.972981 -0.894474 0.7107696 -0.040478 -0.959527 
0.8436530 1.4981862 0.8285582 -1.284187 1.3557655 
-0.104296 0.0008397 1.0366740 -0.560620 0.3317805 
-0.869832 -0.542603 0.0047614 -0.015730 -0.781197 
-0.950503 -1.263876 -0.137503 0.1807592 -1.309778 
-0.344607 -0.274737 -0.974701 -0.388816 -0.404218 
-0.440296 -0.242987 -0.795658 1.0049424 -0.713076 
-0.884549 -1.157423 -0.739342 0.5376579 -1.003894 
0.5845880 1.1563029 1.2341283 -1.112798 1.0263674 
0.3489540 -0.630812 -1.465495 1.5165928 -0.757728 
0.3068344 0.3210119 -0.209924 0.2683466 0.1360334 
0.6842508 0.5776563 0.1792170 -0.410341 0.5257919 
-0.825438 -1.360007 -1.768370 0.6737023 -1.277090 
0.1033852 -0.528836 -0.989316 1.0431975 -0.702090 
-0.488006 -0.446422 -0.634326 -1.014849 -0.496939 
0.4536771 0.7061773 0.5050520 -1.175437 0.6949161 
0.2455717 -1.192096 -1.993114 2.0464056 -1.057809 
0.7345045 0.2895936 -0.980236 0.0326499 0.0871396 
0.8792375 1.1271915 -0.071120 -1.148992 0.9628835 
-0.140260 -1.031195 -0.639683 1.6544627 -1.051562 
0.7902142 0.6874468 -0.280460 0.6193673 0.7991353 
0.1693623 0.2599640 -0.229633 0.2807456 0.0711080 
0.1070385 0.2186336 0.4768717 0.1375966 -0.020256 
-0.570264 0.0227951 0.6424880 -1.613961 -0.079706 

